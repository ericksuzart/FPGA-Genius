// The purpose of this module is to select the appropriate pixel, address, and
// clock signals based on the SELECTOR input. It functions as a demultiplexer
// for memory locations, allowing the selection of a specific memory location
// and retrieving the corresponding data from that location.
module MemoryDemux
(
  input [2:0] SELECTOR,
  input [15:0] IN_ADDR,
  input IN_CLK,

  // ----- Input Pixels -----
  input [15:0] BACKGROUND_PX,
  input [15:0] POWER_BTN_PX,
  input [15:0] RED_BTN_PX,
  input [15:0] GREEN_BTN_PX,
  input [15:0] BLUE_BTN_PX,
  input [15:0] YELLOW_BTN_PX,
  input [15:0] WIN_SCREEN_PX,
  input [15:0] LOSE_SCREEN_PX,

  output reg [15:0] OUT_PX,

  // ----- Adresses -----
  output reg [15:0] BACKGROUND_ADDR,  // MAX = 64800
  output reg [15:0] POWER_BTN_ADDR,   // TODO define the MAX =
  output reg [15:0] RED_BTN_ADDR,     // TODO define the MAX =
  output reg [15:0] GREEN_BTN_ADDR,   // TODO define the MAX =
  output reg [15:0] BLUE_BTN_ADDR,    // TODO define the MAX =
  output reg [15:0] YELLOW_BTN_ADDR,  // TODO define the MAX =
  output reg [15:0] WIN_SCREEN_ADDR,  // TODO define the MAX =
  output reg [15:0] LOSE_SCREEN_ADDR, // TODO define the MAX =

  // ----- Clocks -----
  output reg BACKGROUND_CLK,
  output reg POWER_BTN_CLK,
  output reg RED_BTN_CLK,
  output reg GREEN_BTN_CLK,
  output reg BLUE_BTN_CLK,
  output reg YELLOW_BTN_CLK,
  output reg WIN_SCREEN_CLK,
  output reg LOSE_SCREEN_CLK
);

  parameter   BACKGROUND = 3'b000,
              POWER_BTN_ON = 3'b001,
              RED_BTN_ON = 3'b010,
              GREEN_BTN_ON = 3'b011,
              BLUE_BTN_ON = 3'b100,
              YELLOW_BTN_ON = 3'b101,
              WIN_SCREEN = 3'b110,
              LOSE_SCREEN = 3'b111;

  always @(*)
  begin
    OUT_PX = 0;
    BACKGROUND_ADDR = 0;
    BACKGROUND_CLK = 0;
    POWER_BTN_ADDR = 0;
    POWER_BTN_CLK = 0;
    RED_BTN_ADDR = 0;
    RED_BTN_CLK = 0;
    GREEN_BTN_ADDR = 0;
    GREEN_BTN_CLK = 0;
    BLUE_BTN_ADDR = 0;
    BLUE_BTN_CLK = 0;
    YELLOW_BTN_ADDR = 0;
    YELLOW_BTN_CLK = 0;
    WIN_SCREEN_ADDR = 0;
    WIN_SCREEN_CLK = 0;
    LOSE_SCREEN_ADDR = 0;
    LOSE_SCREEN_CLK = 0;

    case (SELECTOR)
      BACKGROUND:
      begin
        OUT_PX = BACKGROUND_PX;
        BACKGROUND_ADDR = IN_ADDR;
        BACKGROUND_CLK = IN_CLK;
      end

      POWER_BTN_ON:
      begin
        OUT_PX = POWER_BTN_PX;
        POWER_BTN_ADDR = IN_ADDR;
        POWER_BTN_CLK = IN_CLK;
      end

      RED_BTN_ON:
      begin
        OUT_PX = RED_BTN_PX;
        RED_BTN_ADDR = IN_ADDR;
        RED_BTN_CLK = IN_CLK;
      end

      GREEN_BTN_ON:
      begin
        OUT_PX = GREEN_BTN_PX;
        GREEN_BTN_ADDR = IN_ADDR;
        GREEN_BTN_CLK = IN_CLK;
      end

      BLUE_BTN_ON:
      begin
        OUT_PX = BLUE_BTN_PX;
        BLUE_BTN_ADDR = IN_ADDR;
        BLUE_BTN_CLK = IN_CLK;
      end

      YELLOW_BTN_ON:
      begin
        OUT_PX = YELLOW_BTN_PX;
        YELLOW_BTN_ADDR = IN_ADDR;
        YELLOW_BTN_CLK = IN_CLK;
      end

      WIN_SCREEN:
      begin
        OUT_PX = WIN_SCREEN_PX;
        WIN_SCREEN_ADDR = IN_ADDR;
        WIN_SCREEN_CLK = IN_CLK;
      end

      LOSE_SCREEN:
      begin
        OUT_PX = LOSE_SCREEN_PX;
        LOSE_SCREEN_ADDR = IN_ADDR;
        LOSE_SCREEN_CLK = IN_CLK;
      end
    endcase
  end
endmodule
